`timescale 1ns/1ns
`include "Capstone.v"

module accumulator_shift_regTB; //Testbench for accumulator
	
endmodule