module Top (input St, input CLK); // control circuit
	
endmodule


module Accumulator (input Si, input Sh, output Xi);

endmodule

module Addend (input Si, input SH, output Yi); //

endmodule

module FullAdder (input x, input y, input Ci, output Si, output Cout); //full adder with flip flop

endmodule






module testbench;
	
endmodule