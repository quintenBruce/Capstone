`timescale 1ns/1ns
`include "Capstone.v"

module addend_shift_regTB; //Testbench for addend
	
endmodule