module Top (input St, input CLK); // control circuit
	
endmodule


module Accumulator (input Si, input Sh, output Xi); // Accumulator

endmodule

module Addend (input Si, input SH, output Yi); // Addend

endmodule

module FullAdder (input x, input y, input Cin, output Si, output Cout); //full adder with flip flop

endmodule



module TopTb; //testbench for entire circuit
	
endmodule

module AccumulatorTb; //testbench for accumulator
	
endmodule

module AddendTb; //testbench for addend
	
endmodule

module FullAdderTb; //testbench for full adder
	
endmodule